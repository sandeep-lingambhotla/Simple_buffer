interface simple_intf();
  bit clk;
  bit reset;
  bit in;
  bit out;
endinterface
