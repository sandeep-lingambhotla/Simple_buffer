//`include "simple_intf.sv"
//interface simple_intf_hrns();
  
//  simple_intf intf(
//   .clk    (dut.clk),
//    .reset  (dut.reset),
//    .in     (dut.in),
//    .out    (dut.out),
//  );
  
//  initial begin  
//    uvm_config_db #(virtual interface simple_intf)::set(null, "*", "simple_vif", simple_intf);
//  end
      
//endinterface
  
//bind simple simple_intf_hrns u_simple_intf_hrns();
